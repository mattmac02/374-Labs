 module encoder(output reg[4:0] Sout, input[31:0] register);
	always @(register)
	begin
		if(register==32'b00000000000000000000000000000001)Sout=0;
		else if(register==32'b00000000000000000000000000000010)Sout=1;
		else if(register==32'b00000000000000000000000000000100)Sout=2;
		else if(register==32'b00000000000000000000000000001000)Sout=3;
		else if(register==32'b00000000000000000000000000010000)Sout=4;
		else if(register==32'b00000000000000000000000000100000)Sout=5;
		else if(register==32'b00000000000000000000000001000000)Sout=6;
		else if(register==32'b00000000000000000000000010000000)Sout=7;
		else if(register==32'b00000000000000000000000100000000)Sout=8;
		else if(register==32'b00000000000000000000001000000000)Sout=9;
		else if(register==32'b00000000000000000000010000000000)Sout=10;
		else if(register==32'b00000000000000000000100000000000)Sout=11;
		else if(register==32'b00000000000000000001000000000000)Sout=12;
		else if(register==32'b00000000000000000010000000000000)Sout=13;
		else if(register==32'b00000000000000000100000000000000)Sout=14;
		else if(register==32'b00000000000000001000000000000000)Sout=15;
		else if(register==32'b00000000000000010000000000000000)Sout=16;
		else if(register==32'b00000000000000100000000000000000)Sout=17;
		else if(register==32'b00000000000001000000000000000000)Sout=18;
		else if(register==32'b00000000000010000000000000000000)Sout=19;
		else if(register==32'b00000000000100000000000000000000)Sout=20;
		else if(register==32'b00000000001000000000000000000000)Sout=21;
		else if(register==32'b00000000010000000000000000000000)Sout=22;
		else if(register==32'b00000000100000000000000000000000)Sout=23;
		else if(register==32'b00000001000000000000000000000000)Sout=24;
		else if(register==32'b00000010000000000000000000000000)Sout=25;
		else if(register==32'b00000100000000000000000000000000)Sout=26;
		else if(register==32'b00001000000000000000000000000000)Sout=27;
		else if(register==32'b00010000000000000000000000000000)Sout=28;
		else if(register==32'b00100000000000000000000000000000)Sout=29;
		else if(register==32'b01000000000000000000000000000000)Sout=30;
		else if(register==32'b10000000000000000000000000000000)Sout=31; else Sout = 5'bx;
	end 

endmodule
